-- Top level for PPM capture and generation
-- Should instantiate both components and map to regs

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.ppm_package.all;

entity ppm_top is

end ppm_top;

architecture structural of ppm_top is



end structural;